magic
tech $PDK
magscale 1 2
timestamp 1606502073
<< metal3 >>
rect -3136 3072 3136 3100
rect -3136 -3072 3052 3072
rect 3116 -3072 3136 3072
rect -3136 -3100 3136 -3072
<< via3 >>
rect 3052 -3072 3116 3072
<< mimcap >>
rect -3036 2960 2964 3000
rect -3036 -2960 2332 2960
rect 2924 -2960 2964 2960
rect -3036 -3000 2964 -2960
<< mimcapcontact >>
rect 2332 -2960 2924 2960
<< metal4 >>
rect 3036 3072 3132 3088
rect 2331 2960 2925 2961
rect 2331 -2960 2332 2960
rect 2924 -2960 2925 2960
rect 2331 -2961 2925 -2960
rect 3036 -3072 3052 3072
rect 3116 -3072 3132 3072
rect 3036 -3088 3132 -3072
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX -3136 -3100 3064 3100
string parameters w 30.00 l 30.00 val 920.4 carea 1.00 cperi 0.17 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov -10
string library sky130
<< end >>
